// tb_exp_lut_unit.v
`timescale 1ns / 1ps

module tb_exp_lut_unit;

    // Parameters from user's exp_lut_unit.v
    parameter INPUT_WIDTH_TB      = 12;
    parameter INPUT_FRAC_BITS_TB  = 8;  // Q4.8 for x_in (S III . FFFFFFFF)
    parameter OUTPUT_WIDTH_TB     = 16;
    parameter OUTPUT_FRAC_BITS_TB = 15; // Q1.15 for y_out (S . FFFFFFFFFFFFFFF)
    parameter LUT_ADDR_WIDTH_TB   = 8;
    parameter EXP_LUT_LATENCY_TB  = 1;
    
    localparam CLK_PERIOD          = 10;

    // DUT Interface Signals
    reg                               clk_tb;
    reg                               rst_n_tb;
    reg                               start_exp_tb;
    reg signed [INPUT_WIDTH_TB-1:0]   x_in_tb;

    wire [OUTPUT_WIDTH_TB-1:0]        y_out_dut; 
    wire                              exp_done_dut;

    // Instantiate the DUT
    exp_lut_unit #(
        .INPUT_WIDTH(INPUT_WIDTH_TB),
        .INPUT_FRAC_BITS(INPUT_FRAC_BITS_TB),
        .OUTPUT_WIDTH(OUTPUT_WIDTH_TB),
        .OUTPUT_FRAC_BITS(OUTPUT_FRAC_BITS_TB),
        .LUT_ADDR_WIDTH(LUT_ADDR_WIDTH_TB),
        .EXP_LUT_LATENCY(EXP_LUT_LATENCY_TB)
    ) DUT (
        .clk(clk_tb),
        .rst_n(rst_n_tb),
        .start_exp(start_exp_tb),
        .x_in(x_in_tb),
        .y_out(y_out_dut), 
        .exp_done(exp_done_dut)
    );

    // Clock generation
    always #(CLK_PERIOD/2) clk_tb = ~clk_tb;

    // Test sequence
    initial begin
        integer timeout_counter;
        reg [OUTPUT_WIDTH_TB-1:0] expected_y_out; 
        real x_real_val;
        logic test_passed_overall; // Declaration moved to top

        clk_tb = 1'b0;
        rst_n_tb = 1'b0;
        start_exp_tb = 1'b0;
        x_in_tb = 0;
        test_passed_overall = 1'b1; // Initialization after declarations

        $display("[%0t TB] Starting Exp LUT Unit Testbench...", $time);
        $display("[%0t TB] NOTE: This TB assumes exp_lut.mem is generated by your Python script.", $time);
        $display("[%0t TB] And that DUT output y_out is effectively UQ0.15 (unsigned with 15 fractional bits).", $time);


        #(CLK_PERIOD * 2);
        rst_n_tb = 1'b1;
        $display("[%0t TB] Reset de-asserted.", $time);
        #(CLK_PERIOD);

        // --- Test Case 1: x_in = 0.0 ---
        // Python script for i=0: x=0, y=exp(0)=1.0. fixed_val = round(1.0 * (2^15)) = 32768 -> 16'h8000
        // DUT for x_in_r == 0: lut_out_comb = (1 << OUTPUT_FRAC_BITS) = (1 << 15) = 16'h8000
        $display("[%0t TB] === Test Case 1: x_in = 0.0 (Q4.8: 0) ===", $time);
        x_real_val = 0.0;
        x_in_tb = $rtoi(x_real_val * (1 << INPUT_FRAC_BITS_TB)); 
        expected_y_out = 16'h8000; 

        start_exp_tb = 1'b1; @(posedge clk_tb); start_exp_tb = 1'b0;
        timeout_counter = 0;
        while (!exp_done_dut && timeout_counter < (EXP_LUT_LATENCY_TB + 5)) begin @(posedge clk_tb); timeout_counter = timeout_counter + 1; end

        if (!exp_done_dut) $error("TC1 TIMEOUT");
        else if (y_out_dut === expected_y_out) $display("TC1 PASSED. x_in=%d, y_out=%h (Exp: %h)", x_in_tb, y_out_dut, expected_y_out);
        else begin $error("TC1 FAILED. x_in=%d, y_out=%h (Exp: %h)", x_in_tb, y_out_dut, expected_y_out); test_passed_overall = 1'b0; end
        #(CLK_PERIOD * 2);

        // --- Test Case 2: x_in = -1 (Q4.8, real -0.00390625) ---
        // Python script: i=1, x=1/256. y=exp(-1/256) ~ 0.996099. fixed_val = round(0.996099 * 2^15) = 32640 (16'h7F80)
        // DUT: abs_x = 1. integer_part = 0. lut_addr_from_frac_part = 1. lut[1] should be 16'h7F80.
        $display("[%0t TB] === Test Case 2: x_in = -1 (Q4.8, real -0.00390625) ===", $time);
        x_real_val = -1.0/256.0;
        x_in_tb = $rtoi(x_real_val * (1 << INPUT_FRAC_BITS_TB)); 
        expected_y_out = 16'h7F80; // From Python script logic for i=1

        start_exp_tb = 1'b1; @(posedge clk_tb); start_exp_tb = 1'b0;
        timeout_counter = 0;
        while (!exp_done_dut && timeout_counter < (EXP_LUT_LATENCY_TB + 5)) begin @(posedge clk_tb); timeout_counter = timeout_counter + 1; end

        if (!exp_done_dut) $error("TC2 TIMEOUT");
        else if (y_out_dut === expected_y_out) $display("TC2 PASSED. x_in=%d, y_out=%h (Exp: %h)", x_in_tb, y_out_dut, expected_y_out);
        else begin $error("TC2 FAILED. x_in=%d, y_out=%h (Exp: %h)", x_in_tb, y_out_dut, expected_y_out); test_passed_overall = 1'b0; end
        #(CLK_PERIOD * 2);

        // --- Test Case 3: x_in = -128 (Q4.8, real -0.5) ---
        // Python script: i=128, x=128/256=0.5. y=exp(-0.5) ~ 0.60653. fixed_val = round(0.60653 * 2^15) = 19875 (16'h4D9F)
        // DUT: abs_x = 128. integer_part = 0. lut_addr_from_frac_part = 128. lut[128] should be 16'h4D9F.
        $display("[%0t TB] === Test Case 3: x_in = -128 (Q4.8, real -0.5) ===", $time);
        x_real_val = -0.5;
        x_in_tb = $rtoi(x_real_val * (1 << INPUT_FRAC_BITS_TB)); 
        expected_y_out = 16'h4D9F;

        start_exp_tb = 1'b1; @(posedge clk_tb); start_exp_tb = 1'b0;
        timeout_counter = 0;
        while (!exp_done_dut && timeout_counter < (EXP_LUT_LATENCY_TB + 5)) begin @(posedge clk_tb); timeout_counter = timeout_counter + 1; end

        if (!exp_done_dut) $error("TC3 TIMEOUT");
        else if (y_out_dut === expected_y_out) $display("TC3 PASSED. x_in=%d, y_out=%h (Exp: %h)", x_in_tb, y_out_dut, expected_y_out);
        else begin $error("TC3 FAILED. x_in=%d, y_out=%h (Exp: %h)", x_in_tb, y_out_dut, expected_y_out); test_passed_overall = 1'b0; end
        #(CLK_PERIOD * 2);
        
        // --- Test Case 4: x_in very negative (e.g. -2.0) ---
        // Input x_in (Q4.8) = -2.0 * 256 = -512
        // DUT: abs_x = 512. integer_part_of_abs_x = 2 (non-zero).
        // DUT should output OUTPUT_WIDTH'(1) = 16'h0001
        $display("[%0t TB] === Test Case 4: x_in = -2.0 (Q4.8: -512) ===", $time);
        x_real_val = -2.0;
        x_in_tb = $rtoi(x_real_val * (1 << INPUT_FRAC_BITS_TB)); 
        expected_y_out = 16'h0001; 

        start_exp_tb = 1'b1; @(posedge clk_tb); start_exp_tb = 1'b0;
        timeout_counter = 0;
        while (!exp_done_dut && timeout_counter < (EXP_LUT_LATENCY_TB + 5)) begin @(posedge clk_tb); timeout_counter = timeout_counter + 1; end

        if (!exp_done_dut) $error("TC4 TIMEOUT");
        else if (y_out_dut === expected_y_out) $display("TC4 PASSED. x_in=%d, y_out=%h (Exp: %h)", x_in_tb, y_out_dut, expected_y_out);
        else begin $error("TC4 FAILED. x_in=%d, y_out=%h (Exp: %h)", x_in_tb, y_out_dut, expected_y_out); test_passed_overall = 1'b0; end
        #(CLK_PERIOD * 5); 


        if(test_passed_overall) $display("[%0t TB] ALL EXP LUT TEST CASES PASSED.", $time);
        else $display("[%0t TB] ONE OR MORE EXP LUT TEST CASES FAILED.", $time);

        $display("[%0t TB] Exp LUT Unit Testbench Finished.", $time);
        $finish;
    end

endmodule

