// exp_lut_unit.v (Corrected LUT Addressing and Logic for User's Parameters)
module exp_lut_unit #(
    parameter INPUT_WIDTH         = 12, // Q4.8 (S III FFFFFFFF)
    parameter INPUT_FRAC_BITS     = 8,
    parameter OUTPUT_WIDTH        = 16, // Q1.15 (S .FFFFFFFFFFFFFFF) per TB expectation
    parameter OUTPUT_FRAC_BITS    = 15,
    parameter LUT_ADDR_WIDTH      = 8,   // 256 entries, matches Python script's N
    parameter EXP_LUT_LATENCY     = 1
)(
    input  wire                          clk,
    input  wire                          rst_n,
    input  wire                          start_exp,
    input  wire signed [INPUT_WIDTH-1:0] x_in,

    output reg [OUTPUT_WIDTH-1:0]        y_out,    // Matched to user's TB (unsigned)
    output reg                           exp_done
);

    reg signed [INPUT_WIDTH-1:0] x_in_r;
    reg [EXP_LUT_LATENCY:0]      latency_counter_reg;
    reg                          exp_done_pulse_reg;

    wire [INPUT_WIDTH-1:0]     abs_x_comb = (x_in_r[INPUT_WIDTH-1] && x_in_r != 0) ? -x_in_r : x_in_r;
    
    // Integer part of abs_x (e.g., bits [11:8] for Q4.8)
    wire [INPUT_WIDTH-1-INPUT_FRAC_BITS:0] abs_x_integer_part = abs_x_comb[INPUT_WIDTH-1 : INPUT_FRAC_BITS];
    
    // Fractional part of abs_x (e.g., bits [7:0] for Q4.8) used for LUT address
    wire [LUT_ADDR_WIDTH-1:0] lut_addr_calc;
    // Python script uses i from 0 to N-1 (255) as address, where x_for_exp = i / (2^FRAC_BITS)
    // So, if abs_x_comb < 1.0, its fractional part scaled by 2^FRAC_BITS is the address.
    // Since LUT_ADDR_WIDTH == INPUT_FRAC_BITS here, we use all fractional bits.
    assign lut_addr_calc = abs_x_comb[INPUT_FRAC_BITS-1 : 0];


    reg [OUTPUT_WIDTH-1:0] lut [0:(1<<LUT_ADDR_WIDTH)-1];
    initial begin
        $display("[%0t EXP_LUT_DUT] Reading exp_lut.mem (LUT_SIZE=%d)...", $time, (1<<LUT_ADDR_WIDTH));
        $readmemh("exp_lut.mem", lut); // Generated by Python script
    end

    wire [OUTPUT_WIDTH-1:0] lut_out_comb;

    // LUT lookup logic
    assign lut_out_comb = (x_in_r == 0) ? OUTPUT_WIDTH'(1 << OUTPUT_FRAC_BITS) : // exp(0) = 1.0
                        (x_in_r > 0) ? OUTPUT_WIDTH'(1) : // Error/Smallest: Input should be <=0
                        (|abs_x_integer_part) ? OUTPUT_WIDTH'(1) : // If abs(x_in_r) >= 1.0, exp(-abs(x)) is small
                                                                   // Python LUT only covers abs(x) in [0, 1)
                        lut[lut_addr_calc]; // Use fractional part as address if abs(x_in_r) < 1.0

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            x_in_r <= 0;
            y_out <= 0;
            exp_done <= 1'b0;
            latency_counter_reg <= 0;
            exp_done_pulse_reg <= 1'b0;
        end else begin
            exp_done_pulse_reg <= 1'b0;

            if (start_exp) begin
                x_in_r <= x_in;
                if (EXP_LUT_LATENCY == 0) begin
                    y_out <= lut_out_comb;
                    exp_done_pulse_reg <= 1'b1;
                end else begin
                    latency_counter_reg <= EXP_LUT_LATENCY;
                    exp_done <= 1'b0;
                end
            end else if (latency_counter_reg > 0) begin
                latency_counter_reg <= latency_counter_reg - 1;
                if (latency_counter_reg == 1) begin
                    y_out <= lut_out_comb; // lut_out_comb uses x_in_r from start_exp cycle
                    exp_done_pulse_reg <= 1'b1;
                end
            end
            exp_done <= exp_done_pulse_reg;
        end
    end
endmodule

